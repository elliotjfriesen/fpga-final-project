library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
  port(
	  clock : in std_logic;
	  row_count : in unsigned(5 downto 0);
	  col_count : in unsigned(6 downto 0);
	  rgb : out std_logic_vector(5 downto 0)
  );
end rom;

architecture synth of rom is
signal address : unsigned(12 downto 0);
signal rgb_signal : std_logic_vector(5 downto 0);
begin
address <= row_count & col_count;
	process (clock) begin
	if rising_edge(clock) then
rgb_signal <=             "000000" when address = "0001000000101" else
            "000000" when address = "0001000000110" else
            "000000" when address = "0001000000111" else
            "000000" when address = "0001000001100" else
            "000000" when address = "0001000001101" else
            "000000" when address = "0001000001110" else
            "000000" when address = "0001000010011" else
            "000000" when address = "0001000010100" else
            "000000" when address = "0001000011011" else
            "000000" when address = "0001000011100" else
            "000000" when address = "0001000100011" else
            "000000" when address = "0001000100100" else
            "000000" when address = "0001000100101" else
            "000000" when address = "0001000100110" else
            "000000" when address = "0001000100111" else
            "000000" when address = "0001000101000" else
            "000000" when address = "0001000101001" else
            "000000" when address = "0001000101010" else
            "000000" when address = "0001000101111" else
            "000000" when address = "0001000110000" else
            "000000" when address = "0001000110001" else
            "000000" when address = "0001000110010" else
            "000000" when address = "0001000110011" else
            "000000" when address = "0001000110100" else
            "000000" when address = "0001000110101" else
            "000000" when address = "0001000110110" else
            "000000" when address = "0001000111111" else
            "000000" when address = "0001001000000" else
            "000000" when address = "0001001000001" else
            "000000" when address = "0001001000010" else
            "000000" when address = "0001001000011" else
            "000000" when address = "0001001000100" else
            "000000" when address = "0001001000101" else
            "000000" when address = "0001010000101" else
            "000000" when address = "0001010000110" else
            "000000" when address = "0001010000111" else
            "000000" when address = "0001010001000" else
            "000000" when address = "0001010001011" else
            "000000" when address = "0001010001100" else
            "000000" when address = "0001010001101" else
            "000000" when address = "0001010001110" else
            "000000" when address = "0001010010011" else
            "000000" when address = "0001010010100" else
            "000000" when address = "0001010011011" else
            "000000" when address = "0001010011100" else
            "000000" when address = "0001010100010" else
            "000000" when address = "0001010100011" else
            "000000" when address = "0001010100100" else
            "000000" when address = "0001010100101" else
            "000000" when address = "0001010100110" else
            "000000" when address = "0001010100111" else
            "000000" when address = "0001010101000" else
            "000000" when address = "0001010101001" else
            "000000" when address = "0001010101010" else
            "000000" when address = "0001010101111" else
            "000000" when address = "0001010110000" else
            "000000" when address = "0001010110001" else
            "000000" when address = "0001010110010" else
            "000000" when address = "0001010110011" else
            "000000" when address = "0001010110100" else
            "000000" when address = "0001010110101" else
            "000000" when address = "0001010110110" else
            "000000" when address = "0001010111110" else
            "000000" when address = "0001010111111" else
            "000000" when address = "0001011000000" else
            "000000" when address = "0001011000001" else
            "000000" when address = "0001011000010" else
            "000000" when address = "0001011000011" else
            "000000" when address = "0001011000100" else
            "000000" when address = "0001011000101" else
            "000000" when address = "0001100000101" else
            "000000" when address = "0001100000110" else
            "000000" when address = "0001100000111" else
            "000000" when address = "0001100001000" else
            "000000" when address = "0001100001011" else
            "000000" when address = "0001100001100" else
            "000000" when address = "0001100001101" else
            "000000" when address = "0001100001110" else
            "000000" when address = "0001100010011" else
            "000000" when address = "0001100010100" else
            "000000" when address = "0001100011011" else
            "000000" when address = "0001100011100" else
            "000000" when address = "0001100100010" else
            "000000" when address = "0001100100011" else
            "000000" when address = "0001100110010" else
            "000000" when address = "0001100110011" else
            "000000" when address = "0001100111110" else
            "000000" when address = "0001100111111" else
            "000000" when address = "0001110000101" else
            "000000" when address = "0001110000110" else
            "000000" when address = "0001110000111" else
            "000000" when address = "0001110001000" else
            "000000" when address = "0001110001011" else
            "000000" when address = "0001110001100" else
            "000000" when address = "0001110001101" else
            "000000" when address = "0001110001110" else
            "000000" when address = "0001110010011" else
            "000000" when address = "0001110010100" else
            "000000" when address = "0001110011011" else
            "000000" when address = "0001110011100" else
            "000000" when address = "0001110100010" else
            "000000" when address = "0001110100011" else
            "000000" when address = "0001110110010" else
            "000000" when address = "0001110110011" else
            "000000" when address = "0001110111110" else
            "000000" when address = "0001110111111" else
            "000000" when address = "0010000000101" else
            "000000" when address = "0010000000110" else
            "000000" when address = "0010000000111" else
            "000000" when address = "0010000001000" else
            "000000" when address = "0010000001001" else
            "000000" when address = "0010000001010" else
            "000000" when address = "0010000001011" else
            "000000" when address = "0010000001100" else
            "000000" when address = "0010000001101" else
            "000000" when address = "0010000001110" else
            "000000" when address = "0010000010011" else
            "000000" when address = "0010000010100" else
            "000000" when address = "0010000011011" else
            "000000" when address = "0010000011100" else
            "000000" when address = "0010000100010" else
            "000000" when address = "0010000100011" else
            "000000" when address = "0010000100100" else
            "000000" when address = "0010000100101" else
            "000000" when address = "0010000100110" else
            "000000" when address = "0010000100111" else
            "000000" when address = "0010000101000" else
            "000000" when address = "0010000101001" else
            "000000" when address = "0010000110010" else
            "000000" when address = "0010000110011" else
            "000000" when address = "0010000111110" else
            "000000" when address = "0010000111111" else
            "000000" when address = "0010010000101" else
            "000000" when address = "0010010000110" else
            "000000" when address = "0010010001000" else
            "000000" when address = "0010010001001" else
            "000000" when address = "0010010001010" else
            "000000" when address = "0010010001011" else
            "000000" when address = "0010010001101" else
            "000000" when address = "0010010001110" else
            "000000" when address = "0010010010011" else
            "000000" when address = "0010010010100" else
            "000000" when address = "0010010011011" else
            "000000" when address = "0010010011100" else
            "000000" when address = "0010010100011" else
            "000000" when address = "0010010100100" else
            "000000" when address = "0010010100101" else
            "000000" when address = "0010010100110" else
            "000000" when address = "0010010100111" else
            "000000" when address = "0010010101000" else
            "000000" when address = "0010010101001" else
            "000000" when address = "0010010101010" else
            "000000" when address = "0010010110010" else
            "000000" when address = "0010010110011" else
            "000000" when address = "0010010111110" else
            "000000" when address = "0010010111111" else
            "000000" when address = "0010100000101" else
            "000000" when address = "0010100000110" else
            "000000" when address = "0010100001000" else
            "000000" when address = "0010100001001" else
            "000000" when address = "0010100001010" else
            "000000" when address = "0010100001011" else
            "000000" when address = "0010100001101" else
            "000000" when address = "0010100001110" else
            "000000" when address = "0010100010011" else
            "000000" when address = "0010100010100" else
            "000000" when address = "0010100011011" else
            "000000" when address = "0010100011100" else
            "000000" when address = "0010100101001" else
            "000000" when address = "0010100101010" else
            "000000" when address = "0010100110010" else
            "000000" when address = "0010100110011" else
            "000000" when address = "0010100111110" else
            "000000" when address = "0010100111111" else
            "000000" when address = "0010110000101" else
            "000000" when address = "0010110000110" else
            "000000" when address = "0010110001000" else
            "000000" when address = "0010110001001" else
            "000000" when address = "0010110001010" else
            "000000" when address = "0010110001011" else
            "000000" when address = "0010110001101" else
            "000000" when address = "0010110001110" else
            "000000" when address = "0010110010011" else
            "000000" when address = "0010110010100" else
            "000000" when address = "0010110010101" else
            "000000" when address = "0010110011010" else
            "000000" when address = "0010110011011" else
            "000000" when address = "0010110011100" else
            "000000" when address = "0010110101001" else
            "000000" when address = "0010110101010" else
            "000000" when address = "0010110110010" else
            "000000" when address = "0010110110011" else
            "000000" when address = "0010110111110" else
            "000000" when address = "0010110111111" else
            "000000" when address = "0011000000101" else
            "000000" when address = "0011000000110" else
            "000000" when address = "0011000001001" else
            "000000" when address = "0011000001010" else
            "000000" when address = "0011000001101" else
            "000000" when address = "0011000001110" else
            "000000" when address = "0011000010100" else
            "000000" when address = "0011000010101" else
            "000000" when address = "0011000010110" else
            "000000" when address = "0011000010111" else
            "000000" when address = "0011000011000" else
            "000000" when address = "0011000011001" else
            "000000" when address = "0011000011010" else
            "000000" when address = "0011000011011" else
            "000000" when address = "0011000100010" else
            "000000" when address = "0011000100011" else
            "000000" when address = "0011000100100" else
            "000000" when address = "0011000100101" else
            "000000" when address = "0011000100110" else
            "000000" when address = "0011000100111" else
            "000000" when address = "0011000101000" else
            "000000" when address = "0011000101001" else
            "000000" when address = "0011000101010" else
            "000000" when address = "0011000101111" else
            "000000" when address = "0011000110000" else
            "000000" when address = "0011000110001" else
            "000000" when address = "0011000110010" else
            "000000" when address = "0011000110011" else
            "000000" when address = "0011000110100" else
            "000000" when address = "0011000110101" else
            "000000" when address = "0011000110110" else
            "000000" when address = "0011000111110" else
            "000000" when address = "0011000111111" else
            "000000" when address = "0011001000000" else
            "000000" when address = "0011001000001" else
            "000000" when address = "0011001000010" else
            "000000" when address = "0011001000011" else
            "000000" when address = "0011001000100" else
            "000000" when address = "0011001000101" else
            "000000" when address = "0011010000101" else
            "000000" when address = "0011010000110" else
            "000000" when address = "0011010001001" else
            "000000" when address = "0011010001010" else
            "000000" when address = "0011010001101" else
            "000000" when address = "0011010001110" else
            "000000" when address = "0011010010101" else
            "000000" when address = "0011010010110" else
            "000000" when address = "0011010010111" else
            "000000" when address = "0011010011000" else
            "000000" when address = "0011010011001" else
            "000000" when address = "0011010011010" else
            "000000" when address = "0011010100010" else
            "000000" when address = "0011010100011" else
            "000000" when address = "0011010100100" else
            "000000" when address = "0011010100101" else
            "000000" when address = "0011010100110" else
            "000000" when address = "0011010100111" else
            "000000" when address = "0011010101000" else
            "000000" when address = "0011010101001" else
            "000000" when address = "0011010101111" else
            "000000" when address = "0011010110000" else
            "000000" when address = "0011010110001" else
            "000000" when address = "0011010110010" else
            "000000" when address = "0011010110011" else
            "000000" when address = "0011010110100" else
            "000000" when address = "0011010110101" else
            "000000" when address = "0011010110110" else
            "000000" when address = "0011010111111" else
            "000000" when address = "0011011000000" else
            "000000" when address = "0011011000001" else
            "000000" when address = "0011011000010" else
            "000000" when address = "0011011000011" else
            "000000" when address = "0011011000100" else
            "000000" when address = "0011011000101" else
            "000000" when address = "0100110101111" else
            "000000" when address = "0100110110000" else
            "000000" when address = "0100110110001" else
            "000000" when address = "0100110110010" else
            "000000" when address = "0100110110011" else
            "000000" when address = "0100110110100" else
            "000000" when address = "0100110110101" else
            "000000" when address = "0100110111111" else
            "000000" when address = "0100111000000" else
            "000000" when address = "0100111000001" else
            "000000" when address = "0100111000010" else
            "000000" when address = "0100111000011" else
            "000000" when address = "0100111000100" else
            "000000" when address = "0100111000101" else
            "000000" when address = "0101000000101" else
            "000000" when address = "0101000000110" else
            "000000" when address = "0101000000111" else
            "000000" when address = "0101000001000" else
            "000000" when address = "0101000001001" else
            "000000" when address = "0101000001010" else
            "000000" when address = "0101000001011" else
            "000000" when address = "0101000001100" else
            "000000" when address = "0101000001101" else
            "000000" when address = "0101000010100" else
            "000000" when address = "0101000010101" else
            "000000" when address = "0101000010110" else
            "000000" when address = "0101000010111" else
            "000000" when address = "0101000011000" else
            "000000" when address = "0101000011001" else
            "000000" when address = "0101000011010" else
            "000000" when address = "0101000011011" else
            "000000" when address = "0101000100011" else
            "000000" when address = "0101000100100" else
            "000000" when address = "0101000101111" else
            "000000" when address = "0101000110000" else
            "000000" when address = "0101000110001" else
            "000000" when address = "0101000110010" else
            "000000" when address = "0101000110011" else
            "000000" when address = "0101000110100" else
            "000000" when address = "0101000110101" else
            "000000" when address = "0101000111110" else
            "000000" when address = "0101000111111" else
            "000000" when address = "0101001000000" else
            "000000" when address = "0101001000001" else
            "000000" when address = "0101001000010" else
            "000000" when address = "0101001000011" else
            "000000" when address = "0101001000100" else
            "000000" when address = "0101001000101" else
            "000000" when address = "0101010000101" else
            "000000" when address = "0101010000110" else
            "000000" when address = "0101010000111" else
            "000000" when address = "0101010001000" else
            "000000" when address = "0101010001001" else
            "000000" when address = "0101010001010" else
            "000000" when address = "0101010001011" else
            "000000" when address = "0101010001100" else
            "000000" when address = "0101010001101" else
            "000000" when address = "0101010010100" else
            "000000" when address = "0101010010101" else
            "000000" when address = "0101010010110" else
            "000000" when address = "0101010010111" else
            "000000" when address = "0101010011000" else
            "000000" when address = "0101010011001" else
            "000000" when address = "0101010011010" else
            "000000" when address = "0101010011011" else
            "000000" when address = "0101010100011" else
            "000000" when address = "0101010100100" else
            "000000" when address = "0101010101111" else
            "000000" when address = "0101010110000" else
            "000000" when address = "0101010111110" else
            "000000" when address = "0101010111111" else
            "000000" when address = "0101100001001" else
            "000000" when address = "0101100001010" else
            "000000" when address = "0101100010111" else
            "000000" when address = "0101100011000" else
            "000000" when address = "0101100100011" else
            "000000" when address = "0101100100100" else
            "000000" when address = "0101100101111" else
            "000000" when address = "0101100110000" else
            "000000" when address = "0101100111110" else
            "000000" when address = "0101100111111" else
            "000000" when address = "0101110001001" else
            "000000" when address = "0101110001010" else
            "000000" when address = "0101110010111" else
            "000000" when address = "0101110011000" else
            "000000" when address = "0101110100011" else
            "000000" when address = "0101110100100" else
            "000000" when address = "0101110101111" else
            "000000" when address = "0101110110000" else
            "000000" when address = "0101110110001" else
            "000000" when address = "0101110110010" else
            "000000" when address = "0101110110011" else
            "000000" when address = "0101110110100" else
            "000000" when address = "0101110110101" else
            "000000" when address = "0101110111110" else
            "000000" when address = "0101110111111" else
            "000000" when address = "0110000001001" else
            "000000" when address = "0110000001010" else
            "000000" when address = "0110000010111" else
            "000000" when address = "0110000011000" else
            "000000" when address = "0110000100011" else
            "000000" when address = "0110000100100" else
            "000000" when address = "0110000101111" else
            "000000" when address = "0110000110000" else
            "000000" when address = "0110000110001" else
            "000000" when address = "0110000110010" else
            "000000" when address = "0110000110011" else
            "000000" when address = "0110000110100" else
            "000000" when address = "0110000110101" else
            "000000" when address = "0110000111110" else
            "000000" when address = "0110000111111" else
            "000000" when address = "0110001000000" else
            "000000" when address = "0110001000001" else
            "000000" when address = "0110001000010" else
            "000000" when address = "0110001000011" else
            "000000" when address = "0110001000100" else
            "000000" when address = "0110010001001" else
            "000000" when address = "0110010001010" else
            "000000" when address = "0110010010111" else
            "000000" when address = "0110010011000" else
            "000000" when address = "0110010100011" else
            "000000" when address = "0110010100100" else
            "000000" when address = "0110010101111" else
            "000000" when address = "0110010110000" else
            "000000" when address = "0110010111111" else
            "000000" when address = "0110011000000" else
            "000000" when address = "0110011000001" else
            "000000" when address = "0110011000010" else
            "000000" when address = "0110011000011" else
            "000000" when address = "0110011000100" else
            "000000" when address = "0110011000101" else
            "000000" when address = "0110100001001" else
            "000000" when address = "0110100001010" else
            "000000" when address = "0110100010111" else
            "000000" when address = "0110100011000" else
            "000000" when address = "0110100100011" else
            "000000" when address = "0110100100100" else
            "000000" when address = "0110100101111" else
            "000000" when address = "0110100110000" else
            "000000" when address = "0110101000100" else
            "000000" when address = "0110101000101" else
            "000000" when address = "0110110001001" else
            "000000" when address = "0110110001010" else
            "000000" when address = "0110110010111" else
            "000000" when address = "0110110011000" else
            "000000" when address = "0110110100011" else
            "000000" when address = "0110110100100" else
            "000000" when address = "0110110101111" else
            "000000" when address = "0110110110000" else
            "000000" when address = "0110111000100" else
            "000000" when address = "0110111000101" else
            "000000" when address = "0111000001001" else
            "000000" when address = "0111000001010" else
            "000000" when address = "0111000010100" else
            "000000" when address = "0111000010101" else
            "000000" when address = "0111000010110" else
            "000000" when address = "0111000010111" else
            "000000" when address = "0111000011000" else
            "000000" when address = "0111000011001" else
            "000000" when address = "0111000011010" else
            "000000" when address = "0111000011011" else
            "000000" when address = "0111000100011" else
            "000000" when address = "0111000100100" else
            "000000" when address = "0111000100101" else
            "000000" when address = "0111000100110" else
            "000000" when address = "0111000100111" else
            "000000" when address = "0111000101000" else
            "000000" when address = "0111000101001" else
            "000000" when address = "0111000101111" else
            "000000" when address = "0111000110000" else
            "000000" when address = "0111000110001" else
            "000000" when address = "0111000110010" else
            "000000" when address = "0111000110011" else
            "000000" when address = "0111000110100" else
            "000000" when address = "0111000110101" else
            "000000" when address = "0111000111110" else
            "000000" when address = "0111000111111" else
            "000000" when address = "0111001000000" else
            "000000" when address = "0111001000001" else
            "000000" when address = "0111001000010" else
            "000000" when address = "0111001000011" else
            "000000" when address = "0111001000100" else
            "000000" when address = "0111001000101" else
            "000000" when address = "0111010001001" else
            "000000" when address = "0111010001010" else
            "000000" when address = "0111010010100" else
            "000000" when address = "0111010010101" else
            "000000" when address = "0111010010110" else
            "000000" when address = "0111010010111" else
            "000000" when address = "0111010011000" else
            "000000" when address = "0111010011001" else
            "000000" when address = "0111010011010" else
            "000000" when address = "0111010011011" else
            "000000" when address = "0111010100011" else
            "000000" when address = "0111010100100" else
            "000000" when address = "0111010100101" else
            "000000" when address = "0111010100110" else
            "000000" when address = "0111010100111" else
            "000000" when address = "0111010101000" else
            "000000" when address = "0111010101001" else
            "000000" when address = "0111010101111" else
            "000000" when address = "0111010110000" else
            "000000" when address = "0111010110001" else
            "000000" when address = "0111010110010" else
            "000000" when address = "0111010110011" else
            "000000" when address = "0111010110100" else
            "000000" when address = "0111010110101" else
            "000000" when address = "0111010111110" else
            "000000" when address = "0111010111111" else
            "000000" when address = "0111011000000" else
            "000000" when address = "0111011000001" else
            "000000" when address = "0111011000010" else
            "000000" when address = "0111011000011" else
            "000000" when address = "0111011000100" else
            "000000" when address = "1011000000000" else
            "000000" when address = "1011000000001" else
            "000000" when address = "1011000000010" else
            "000000" when address = "1011000000011" else
            "000000" when address = "1011000000100" else
            "000000" when address = "1011000000101" else
            "000000" when address = "1011000000110" else
            "000000" when address = "1011000000111" else
            "000000" when address = "1011000001000" else
            "000000" when address = "1011000001001" else
            "000000" when address = "1011000001010" else
            "000000" when address = "1011000001011" else
            "000000" when address = "1011000001100" else
            "000000" when address = "1011000001101" else
            "000000" when address = "1011000001110" else
            "000000" when address = "1011000001111" else
            "000000" when address = "1011000010000" else
            "000000" when address = "1011000010001" else
            "000000" when address = "1011000010010" else
            "000000" when address = "1011000010011" else
            "000000" when address = "1011000010100" else
            "000000" when address = "1011000010101" else
            "000000" when address = "1011000010110" else
            "000000" when address = "1011000010111" else
            "000000" when address = "1011000011000" else
            "000000" when address = "1011000011001" else
            "000000" when address = "1011000011010" else
            "000000" when address = "1011000011011" else
            "000000" when address = "1011000011100" else
            "000000" when address = "1011000011101" else
            "000000" when address = "1011000011110" else
            "000000" when address = "1011000011111" else
            "000000" when address = "1011000100000" else
            "000000" when address = "1011000100001" else
            "000000" when address = "1011000100010" else
            "000000" when address = "1011000100011" else
            "000000" when address = "1011000100100" else
            "000000" when address = "1011000100101" else
            "000000" when address = "1011000100110" else
            "000000" when address = "1011000100111" else
            "000000" when address = "1011000101000" else
            "000000" when address = "1011000101001" else
            "000000" when address = "1011000101010" else
            "000000" when address = "1011000101011" else
            "000000" when address = "1011000101100" else
            "000000" when address = "1011000101101" else
            "000000" when address = "1011000101110" else
            "000000" when address = "1011000101111" else
            "000000" when address = "1011000110000" else
            "000000" when address = "1011000110001" else
            "000000" when address = "1011000110010" else
            "000000" when address = "1011000110011" else
            "000000" when address = "1011000110100" else
            "000000" when address = "1011000110101" else
            "000000" when address = "1011000110110" else
            "000000" when address = "1011000110111" else
            "000000" when address = "1011000111000" else
            "000000" when address = "1011000111001" else
            "000000" when address = "1011000111010" else
            "000000" when address = "1011000111011" else
            "000000" when address = "1011000111100" else
            "000000" when address = "1011000111101" else
            "000000" when address = "1011000111110" else
            "000000" when address = "1011000111111" else
            "000000" when address = "1011001000000" else
            "000000" when address = "1011001000001" else
            "000000" when address = "1011001000010" else
            "000000" when address = "1011001000011" else
            "000000" when address = "1011001000100" else
            "000000" when address = "1011001000101" else
            "000000" when address = "1011001000110" else
            "000000" when address = "1011001000111" else
            "000000" when address = "1011001001000" else
            "000000" when address = "1011001001001" else
            "000000" when address = "1011001001010" else
            "000000" when address = "1011001001011" else
            "000000" when address = "1011001001100" else
            "000000" when address = "1011001001101" else
            "000000" when address = "1011001001110" else
            "000000" when address = "1011001001111" else
            "000000" when address = "1011010000000" else
            "000000" when address = "1011010000001" else
            "000000" when address = "1011010000010" else
            "000000" when address = "1011010000011" else
            "000000" when address = "1011010000100" else
            "000000" when address = "1011010000101" else
            "000000" when address = "1011010000110" else
            "000000" when address = "1011010000111" else
            "000000" when address = "1011010001000" else
            "000000" when address = "1011010001001" else
            "000000" when address = "1011010001010" else
            "000000" when address = "1011010001011" else
            "000000" when address = "1011010001100" else
            "000000" when address = "1011010001101" else
            "000000" when address = "1011010001110" else
            "000000" when address = "1011010001111" else
            "000000" when address = "1011010010000" else
            "000000" when address = "1011010010001" else
            "000000" when address = "1011010010010" else
            "000000" when address = "1011010010011" else
            "000000" when address = "1011010010100" else
            "000000" when address = "1011010010101" else
            "000000" when address = "1011010010110" else
            "000000" when address = "1011010010111" else
            "000000" when address = "1011010011000" else
            "000000" when address = "1011010011001" else
            "000000" when address = "1011010011010" else
            "000000" when address = "1011010011011" else
            "000000" when address = "1011010011100" else
            "000000" when address = "1011010011101" else
            "000000" when address = "1011010011110" else
            "000000" when address = "1011010011111" else
            "000000" when address = "1011010100000" else
            "000000" when address = "1011010100001" else
            "000000" when address = "1011010100010" else
            "000000" when address = "1011010100011" else
            "000000" when address = "1011010100100" else
            "000000" when address = "1011010100101" else
            "000000" when address = "1011010100110" else
            "000000" when address = "1011010100111" else
            "000000" when address = "1011010101000" else
            "000000" when address = "1011010101001" else
            "000000" when address = "1011010101010" else
            "000000" when address = "1011010101011" else
            "000000" when address = "1011010101100" else
            "000000" when address = "1011010101101" else
            "000000" when address = "1011010101110" else
            "000000" when address = "1011010101111" else
            "000000" when address = "1011010110000" else
            "000000" when address = "1011010110001" else
            "000000" when address = "1011010110010" else
            "000000" when address = "1011010110011" else
            "000000" when address = "1011010110100" else
            "000000" when address = "1011010110101" else
            "000000" when address = "1011010110110" else
            "000000" when address = "1011010110111" else
            "000000" when address = "1011010111000" else
            "000000" when address = "1011010111001" else
            "000000" when address = "1011010111010" else
            "000000" when address = "1011010111011" else
            "000000" when address = "1011010111100" else
            "000000" when address = "1011010111101" else
            "000000" when address = "1011010111110" else
            "000000" when address = "1011010111111" else
            "000000" when address = "1011011000000" else
            "000000" when address = "1011011000001" else
            "000000" when address = "1011011000010" else
            "000000" when address = "1011011000011" else
            "000000" when address = "1011011000100" else
            "000000" when address = "1011011000101" else
            "000000" when address = "1011011000110" else
            "000000" when address = "1011011000111" else
            "000000" when address = "1011011001000" else
            "000000" when address = "1011011001001" else
            "000000" when address = "1011011001010" else
            "000000" when address = "1011011001011" else
            "000000" when address = "1011011001100" else
            "000000" when address = "1011011001101" else
            "000000" when address = "1011011001110" else
            "000000" when address = "1011011001111" else
            "000000" when address = "1011100000111" else
            "000000" when address = "1011100001000" else
            "000000" when address = "1011100001001" else
            "000000" when address = "1011100001010" else
            "000000" when address = "1011100010001" else
            "000000" when address = "1011100010010" else
            "000000" when address = "1011100010011" else
            "000000" when address = "1011100010100" else
            "000000" when address = "1011100011011" else
            "000000" when address = "1011100011100" else
            "000000" when address = "1011100011101" else
            "000000" when address = "1011100011110" else
            "000000" when address = "1011100100101" else
            "000000" when address = "1011100100110" else
            "000000" when address = "1011100100111" else
            "000000" when address = "1011100101000" else
            "000000" when address = "1011100101111" else
            "000000" when address = "1011100110000" else
            "000000" when address = "1011100110001" else
            "000000" when address = "1011100110010" else
            "000000" when address = "1011100111001" else
            "000000" when address = "1011100111010" else
            "000000" when address = "1011100111011" else
            "000000" when address = "1011100111100" else
            "000000" when address = "1011101000100" else
            "000000" when address = "1011101000101" else
            "000000" when address = "1011101000110" else
            "000000" when address = "1011101000111" else
            "000000" when address = "1011110000111" else
            "000000" when address = "1011110001000" else
            "000000" when address = "1011110001001" else
            "000000" when address = "1011110001010" else
            "000000" when address = "1011110010001" else
            "000000" when address = "1011110010010" else
            "000000" when address = "1011110010011" else
            "000000" when address = "1011110010100" else
            "000000" when address = "1011110011011" else
            "000000" when address = "1011110011100" else
            "000000" when address = "1011110011101" else
            "000000" when address = "1011110011110" else
            "000000" when address = "1011110100101" else
            "000000" when address = "1011110100110" else
            "000000" when address = "1011110100111" else
            "000000" when address = "1011110101000" else
            "000000" when address = "1011110101111" else
            "000000" when address = "1011110110000" else
            "000000" when address = "1011110110001" else
            "000000" when address = "1011110110010" else
            "000000" when address = "1011110111001" else
            "000000" when address = "1011110111010" else
            "000000" when address = "1011110111011" else
            "000000" when address = "1011110111100" else
            "000000" when address = "1011111000100" else
            "000000" when address = "1011111000101" else
            "000000" when address = "1011111000110" else
            "000000" when address = "1011111000111" else
            "000000" when address = "1100000000111" else
            "000000" when address = "1100000001000" else
            "000000" when address = "1100000001001" else
            "000000" when address = "1100000001010" else
            "000000" when address = "1100000010001" else
            "000000" when address = "1100000010010" else
            "000000" when address = "1100000010011" else
            "000000" when address = "1100000010100" else
            "000000" when address = "1100000011011" else
            "000000" when address = "1100000011100" else
            "000000" when address = "1100000011101" else
            "000000" when address = "1100000011110" else
            "000000" when address = "1100000100101" else
            "000000" when address = "1100000100110" else
            "000000" when address = "1100000100111" else
            "000000" when address = "1100000101000" else
            "000000" when address = "1100000101111" else
            "000000" when address = "1100000110000" else
            "000000" when address = "1100000110001" else
            "000000" when address = "1100000110010" else
            "000000" when address = "1100000111001" else
            "000000" when address = "1100000111010" else
            "000000" when address = "1100000111011" else
            "000000" when address = "1100000111100" else
            "000000" when address = "1100001000100" else
            "000000" when address = "1100001000101" else
            "000000" when address = "1100001000110" else
            "000000" when address = "1100001000111" else
            "000000" when address = "1100010000111" else
            "000000" when address = "1100010001000" else
            "000000" when address = "1100010001001" else
            "000000" when address = "1100010001010" else
            "000000" when address = "1100010010001" else
            "000000" when address = "1100010010010" else
            "000000" when address = "1100010010011" else
            "000000" when address = "1100010010100" else
            "000000" when address = "1100010011011" else
            "000000" when address = "1100010011100" else
            "000000" when address = "1100010011101" else
            "000000" when address = "1100010011110" else
            "000000" when address = "1100010100101" else
            "000000" when address = "1100010100110" else
            "000000" when address = "1100010100111" else
            "000000" when address = "1100010101000" else
            "000000" when address = "1100010101111" else
            "000000" when address = "1100010110000" else
            "000000" when address = "1100010110001" else
            "000000" when address = "1100010110010" else
            "000000" when address = "1100010111001" else
            "000000" when address = "1100010111010" else
            "000000" when address = "1100010111011" else
            "000000" when address = "1100010111100" else
            "000000" when address = "1100011000100" else
            "000000" when address = "1100011000101" else
            "000000" when address = "1100011000110" else
            "000000" when address = "1100011000111" else
            "000000" when address = "1100100000111" else
            "000000" when address = "1100100001000" else
            "000000" when address = "1100100001001" else
            "000000" when address = "1100100001010" else
            "000000" when address = "1100100010001" else
            "000000" when address = "1100100010010" else
            "000000" when address = "1100100010011" else
            "000000" when address = "1100100010100" else
            "000000" when address = "1100100011011" else
            "000000" when address = "1100100011100" else
            "000000" when address = "1100100011101" else
            "000000" when address = "1100100011110" else
            "000000" when address = "1100100100101" else
            "000000" when address = "1100100100110" else
            "000000" when address = "1100100100111" else
            "000000" when address = "1100100101000" else
            "000000" when address = "1100100101111" else
            "000000" when address = "1100100110000" else
            "000000" when address = "1100100110001" else
            "000000" when address = "1100100110010" else
            "000000" when address = "1100100111001" else
            "000000" when address = "1100100111010" else
            "000000" when address = "1100100111011" else
            "000000" when address = "1100100111100" else
            "000000" when address = "1100101000100" else
            "000000" when address = "1100101000101" else
            "000000" when address = "1100101000110" else
            "000000" when address = "1100101000111" else
            "000000" when address = "1100110000111" else
            "000000" when address = "1100110001000" else
            "000000" when address = "1100110001001" else
            "000000" when address = "1100110001010" else
            "000000" when address = "1100110010001" else
            "000000" when address = "1100110010010" else
            "000000" when address = "1100110010011" else
            "000000" when address = "1100110010100" else
            "000000" when address = "1100110011011" else
            "000000" when address = "1100110011100" else
            "000000" when address = "1100110011101" else
            "000000" when address = "1100110011110" else
            "000000" when address = "1100110100101" else
            "000000" when address = "1100110100110" else
            "000000" when address = "1100110100111" else
            "000000" when address = "1100110101000" else
            "000000" when address = "1100110101111" else
            "000000" when address = "1100110110000" else
            "000000" when address = "1100110110001" else
            "000000" when address = "1100110110010" else
            "000000" when address = "1100110111001" else
            "000000" when address = "1100110111010" else
            "000000" when address = "1100110111011" else
            "000000" when address = "1100110111100" else
            "000000" when address = "1100111000100" else
            "000000" when address = "1100111000101" else
            "000000" when address = "1100111000110" else
            "000000" when address = "1100111000111" else
            "000000" when address = "1101000001000" else
            "000000" when address = "1101000001001" else
            "000000" when address = "1101000010010" else
            "000000" when address = "1101000010011" else
            "000000" when address = "1101000011100" else
            "000000" when address = "1101000011101" else
            "000000" when address = "1101000100110" else
            "000000" when address = "1101000100111" else
            "000000" when address = "1101000110000" else
            "000000" when address = "1101000110001" else
            "000000" when address = "1101000111010" else
            "000000" when address = "1101000111011" else
            "000000" when address = "1101001000101" else
            "000000" when address = "1101001000110" else
            "000000" when address = "1101010001000" else
            "000000" when address = "1101010001001" else
            "000000" when address = "1101010010010" else
            "000000" when address = "1101010010011" else
            "000000" when address = "1101010011100" else
            "000000" when address = "1101010011101" else
            "000000" when address = "1101010100110" else
            "000000" when address = "1101010100111" else
            "000000" when address = "1101010110000" else
            "000000" when address = "1101010110001" else
            "000000" when address = "1101010111010" else
            "000000" when address = "1101010111011" else
            "000000" when address = "1101011000101" else
            "000000" when address = "1101011000110" else
            "000000" when address = "1101100001000" else
            "000000" when address = "1101100001001" else
            "000000" when address = "1101100010010" else
            "000000" when address = "1101100010011" else
            "000000" when address = "1101100011100" else
            "000000" when address = "1101100011101" else
            "000000" when address = "1101100100110" else
            "000000" when address = "1101100100111" else
            "000000" when address = "1101100110000" else
            "000000" when address = "1101100110001" else
            "000000" when address = "1101100111010" else
            "000000" when address = "1101100111011" else
            "000000" when address = "1101101000101" else
            "000000" when address = "1101101000110" else
            "000000" when address = "1101110001000" else
            "000000" when address = "1101110001001" else
            "000000" when address = "1101110010010" else
            "000000" when address = "1101110010011" else
            "000000" when address = "1101110011100" else
            "000000" when address = "1101110011101" else
            "000000" when address = "1101110100110" else
            "000000" when address = "1101110100111" else
            "000000" when address = "1101110110000" else
            "000000" when address = "1101110110001" else
            "000000" when address = "1101110111010" else
            "000000" when address = "1101110111011" else
            "000000" when address = "1101111000101" else
            "000000" when address = "1101111000110" else
            "000000" when address = "1110000001000" else
            "000000" when address = "1110000001001" else
            "000000" when address = "1110000010010" else
            "000000" when address = "1110000010011" else
            "000000" when address = "1110000011100" else
            "000000" when address = "1110000011101" else
            "000000" when address = "1110000100110" else
            "000000" when address = "1110000100111" else
            "000000" when address = "1110000110000" else
            "000000" when address = "1110000110001" else
            "000000" when address = "1110000111010" else
            "000000" when address = "1110000111011" else
            "000000" when address = "1110001000101" else
            "000000" when address = "1110001000110" else
            "000000" when address = "1110010001000" else
            "000000" when address = "1110010001001" else
            "000000" when address = "1110010010010" else
            "000000" when address = "1110010010011" else
            "000000" when address = "1110010011100" else
            "000000" when address = "1110010011101" else
            "000000" when address = "1110010100110" else
            "000000" when address = "1110010100111" else
            "000000" when address = "1110010110000" else
            "000000" when address = "1110010110001" else
            "000000" when address = "1110010111010" else
            "000000" when address = "1110010111011" else
            "000000" when address = "1110011000101" else
            "000000" when address = "1110011000110" else
            "000000" when address = "1110100001000" else
            "000000" when address = "1110100001001" else
            "000000" when address = "1110100010010" else
            "000000" when address = "1110100010011" else
            "000000" when address = "1110100011100" else
            "000000" when address = "1110100011101" else
            "000000" when address = "1110100100110" else
            "000000" when address = "1110100100111" else
            "000000" when address = "1110100110000" else
            "000000" when address = "1110100110001" else
            "000000" when address = "1110100111010" else
            "000000" when address = "1110100111011" else
            "000000" when address = "1110101000101" else
            "000000" when address = "1110101000110" else
            "000000" when address = "1110110001000" else
            "000000" when address = "1110110001001" else
            "000000" when address = "1110110010010" else
            "000000" when address = "1110110010011" else
            "000000" when address = "1110110011100" else
            "000000" when address = "1110110011101" else
            "000000" when address = "1110110100110" else
            "000000" when address = "1110110100111" else
            "000000" when address = "1110110110000" else
            "000000" when address = "1110110110001" else
            "000000" when address = "1110110111010" else
            "000000" when address = "1110110111011" else
            "000000" when address = "1110111000101" else
            "000000" when address = "1110111000110" else
                    "111111";



	end if;

	end process;
	
rgb <= rgb_signal;	
			
end;