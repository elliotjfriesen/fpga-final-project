library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gameover is
  port(
	  clock : in std_logic;
	  row_count : in unsigned(5 downto 0);
	  col_count : in unsigned(6 downto 0);
	  rgb : out std_logic_vector(5 downto 0)
  );
end gameover;

architecture synth of gameover is
signal address : unsigned(12 downto 0);
signal rgb_signal : std_logic_vector(5 downto 0);
begin
address <= row_count & col_count;
	process (clock) begin
	if rising_edge(clock) then
rgb_signal <=             "111111" when address = "0000110001101" else
            "111111" when address = "0000110001110" else
            "111111" when address = "0000110001111" else
            "111111" when address = "0000110010000" else
            "111111" when address = "0000110010001" else
            "111111" when address = "0000110010010" else
            "111111" when address = "0000110010011" else
            "111111" when address = "0000110010100" else
            "111111" when address = "0000110011100" else
            "111111" when address = "0000110011101" else
            "111111" when address = "0000110011110" else
            "111111" when address = "0000110011111" else
            "111111" when address = "0000110100000" else
            "111111" when address = "0000110100001" else
            "111111" when address = "0000110101000" else
            "111111" when address = "0000110101001" else
            "111111" when address = "0000110101010" else
            "111111" when address = "0000110110100" else
            "111111" when address = "0000110110101" else
            "111111" when address = "0000110110110" else
            "111111" when address = "0000110111010" else
            "111111" when address = "0000110111011" else
            "111111" when address = "0000110111100" else
            "111111" when address = "0000110111101" else
            "111111" when address = "0000110111110" else
            "111111" when address = "0000110111111" else
            "111111" when address = "0000111000000" else
            "111111" when address = "0000111000001" else
            "111111" when address = "0000111000010" else
            "111111" when address = "0000111000011" else
            "111111" when address = "0000111000100" else
            "111111" when address = "0000111000101" else
            "111111" when address = "0001000001101" else
            "111111" when address = "0001000001110" else
            "111111" when address = "0001000001111" else
            "111111" when address = "0001000010000" else
            "111111" when address = "0001000010001" else
            "111111" when address = "0001000010010" else
            "111111" when address = "0001000010011" else
            "111111" when address = "0001000010100" else
            "111111" when address = "0001000011100" else
            "111111" when address = "0001000011101" else
            "111111" when address = "0001000011110" else
            "111111" when address = "0001000011111" else
            "111111" when address = "0001000100000" else
            "111111" when address = "0001000100001" else
            "111111" when address = "0001000101000" else
            "111111" when address = "0001000101001" else
            "111111" when address = "0001000101010" else
            "111111" when address = "0001000110100" else
            "111111" when address = "0001000110101" else
            "111111" when address = "0001000110110" else
            "111111" when address = "0001000111010" else
            "111111" when address = "0001000111011" else
            "111111" when address = "0001000111100" else
            "111111" when address = "0001000111101" else
            "111111" when address = "0001000111110" else
            "111111" when address = "0001000111111" else
            "111111" when address = "0001001000000" else
            "111111" when address = "0001001000001" else
            "111111" when address = "0001001000010" else
            "111111" when address = "0001001000011" else
            "111111" when address = "0001001000100" else
            "111111" when address = "0001001000101" else
            "111111" when address = "0001010001101" else
            "111111" when address = "0001010001110" else
            "111111" when address = "0001010001111" else
            "111111" when address = "0001010010000" else
            "111111" when address = "0001010010001" else
            "111111" when address = "0001010010010" else
            "111111" when address = "0001010010011" else
            "111111" when address = "0001010010100" else
            "111111" when address = "0001010011100" else
            "111111" when address = "0001010011101" else
            "111111" when address = "0001010011110" else
            "111111" when address = "0001010011111" else
            "111111" when address = "0001010100000" else
            "111111" when address = "0001010100001" else
            "111111" when address = "0001010101000" else
            "111111" when address = "0001010101001" else
            "111111" when address = "0001010101010" else
            "111111" when address = "0001010110100" else
            "111111" when address = "0001010110101" else
            "111111" when address = "0001010110110" else
            "111111" when address = "0001010111010" else
            "111111" when address = "0001010111011" else
            "111111" when address = "0001010111100" else
            "111111" when address = "0001010111101" else
            "111111" when address = "0001010111110" else
            "111111" when address = "0001010111111" else
            "111111" when address = "0001011000000" else
            "111111" when address = "0001011000001" else
            "111111" when address = "0001011000010" else
            "111111" when address = "0001011000011" else
            "111111" when address = "0001011000100" else
            "111111" when address = "0001011000101" else
            "111111" when address = "0001100001010" else
            "111111" when address = "0001100001011" else
            "111111" when address = "0001100001100" else
            "111111" when address = "0001100011001" else
            "111111" when address = "0001100011010" else
            "111111" when address = "0001100011011" else
            "111111" when address = "0001100100010" else
            "111111" when address = "0001100100011" else
            "111111" when address = "0001100100100" else
            "111111" when address = "0001100101000" else
            "111111" when address = "0001100101001" else
            "111111" when address = "0001100101010" else
            "111111" when address = "0001100101011" else
            "111111" when address = "0001100101100" else
            "111111" when address = "0001100101101" else
            "111111" when address = "0001100110001" else
            "111111" when address = "0001100110010" else
            "111111" when address = "0001100110011" else
            "111111" when address = "0001100110100" else
            "111111" when address = "0001100110101" else
            "111111" when address = "0001100110110" else
            "111111" when address = "0001100111010" else
            "111111" when address = "0001100111011" else
            "111111" when address = "0001100111100" else
            "111111" when address = "0001110001010" else
            "111111" when address = "0001110001011" else
            "111111" when address = "0001110001100" else
            "111111" when address = "0001110011001" else
            "111111" when address = "0001110011010" else
            "111111" when address = "0001110011011" else
            "111111" when address = "0001110100010" else
            "111111" when address = "0001110100011" else
            "111111" when address = "0001110100100" else
            "111111" when address = "0001110101000" else
            "111111" when address = "0001110101001" else
            "111111" when address = "0001110101010" else
            "111111" when address = "0001110101011" else
            "111111" when address = "0001110101100" else
            "111111" when address = "0001110101101" else
            "111111" when address = "0001110110001" else
            "111111" when address = "0001110110010" else
            "111111" when address = "0001110110011" else
            "111111" when address = "0001110110100" else
            "111111" when address = "0001110110101" else
            "111111" when address = "0001110110110" else
            "111111" when address = "0001110111010" else
            "111111" when address = "0001110111011" else
            "111111" when address = "0001110111100" else
            "111111" when address = "0010000001010" else
            "111111" when address = "0010000001011" else
            "111111" when address = "0010000001100" else
            "111111" when address = "0010000011001" else
            "111111" when address = "0010000011010" else
            "111111" when address = "0010000011011" else
            "111111" when address = "0010000100010" else
            "111111" when address = "0010000100011" else
            "111111" when address = "0010000100100" else
            "111111" when address = "0010000101000" else
            "111111" when address = "0010000101001" else
            "111111" when address = "0010000101010" else
            "111111" when address = "0010000101011" else
            "111111" when address = "0010000101100" else
            "111111" when address = "0010000101101" else
            "111111" when address = "0010000110001" else
            "111111" when address = "0010000110010" else
            "111111" when address = "0010000110011" else
            "111111" when address = "0010000110100" else
            "111111" when address = "0010000110101" else
            "111111" when address = "0010000110110" else
            "111111" when address = "0010000111010" else
            "111111" when address = "0010000111011" else
            "111111" when address = "0010000111100" else
            "111111" when address = "0010010001010" else
            "111111" when address = "0010010001011" else
            "111111" when address = "0010010001100" else
            "111111" when address = "0010010010000" else
            "111111" when address = "0010010010001" else
            "111111" when address = "0010010010010" else
            "111111" when address = "0010010010011" else
            "111111" when address = "0010010010100" else
            "111111" when address = "0010010010101" else
            "111111" when address = "0010010011001" else
            "111111" when address = "0010010011010" else
            "111111" when address = "0010010011011" else
            "111111" when address = "0010010011100" else
            "111111" when address = "0010010011101" else
            "111111" when address = "0010010011110" else
            "111111" when address = "0010010011111" else
            "111111" when address = "0010010100000" else
            "111111" when address = "0010010100001" else
            "111111" when address = "0010010100010" else
            "111111" when address = "0010010100011" else
            "111111" when address = "0010010100100" else
            "111111" when address = "0010010101000" else
            "111111" when address = "0010010101001" else
            "111111" when address = "0010010101010" else
            "111111" when address = "0010010101110" else
            "111111" when address = "0010010101111" else
            "111111" when address = "0010010110000" else
            "111111" when address = "0010010110100" else
            "111111" when address = "0010010110101" else
            "111111" when address = "0010010110110" else
            "111111" when address = "0010010111010" else
            "111111" when address = "0010010111011" else
            "111111" when address = "0010010111100" else
            "111111" when address = "0010010111101" else
            "111111" when address = "0010010111110" else
            "111111" when address = "0010010111111" else
            "111111" when address = "0010011000000" else
            "111111" when address = "0010011000001" else
            "111111" when address = "0010011000010" else
            "111111" when address = "0010100001010" else
            "111111" when address = "0010100001011" else
            "111111" when address = "0010100001100" else
            "111111" when address = "0010100010000" else
            "111111" when address = "0010100010001" else
            "111111" when address = "0010100010010" else
            "111111" when address = "0010100010011" else
            "111111" when address = "0010100010100" else
            "111111" when address = "0010100010101" else
            "111111" when address = "0010100011001" else
            "111111" when address = "0010100011010" else
            "111111" when address = "0010100011011" else
            "111111" when address = "0010100011100" else
            "111111" when address = "0010100011101" else
            "111111" when address = "0010100011110" else
            "111111" when address = "0010100011111" else
            "111111" when address = "0010100100000" else
            "111111" when address = "0010100100001" else
            "111111" when address = "0010100100010" else
            "111111" when address = "0010100100011" else
            "111111" when address = "0010100100100" else
            "111111" when address = "0010100101000" else
            "111111" when address = "0010100101001" else
            "111111" when address = "0010100101010" else
            "111111" when address = "0010100101110" else
            "111111" when address = "0010100101111" else
            "111111" when address = "0010100110000" else
            "111111" when address = "0010100110100" else
            "111111" when address = "0010100110101" else
            "111111" when address = "0010100110110" else
            "111111" when address = "0010100111010" else
            "111111" when address = "0010100111011" else
            "111111" when address = "0010100111100" else
            "111111" when address = "0010100111101" else
            "111111" when address = "0010100111110" else
            "111111" when address = "0010100111111" else
            "111111" when address = "0010101000000" else
            "111111" when address = "0010101000001" else
            "111111" when address = "0010101000010" else
            "111111" when address = "0010110001010" else
            "111111" when address = "0010110001011" else
            "111111" when address = "0010110001100" else
            "111111" when address = "0010110010000" else
            "111111" when address = "0010110010001" else
            "111111" when address = "0010110010010" else
            "111111" when address = "0010110010011" else
            "111111" when address = "0010110010100" else
            "111111" when address = "0010110010101" else
            "111111" when address = "0010110011001" else
            "111111" when address = "0010110011010" else
            "111111" when address = "0010110011011" else
            "111111" when address = "0010110011100" else
            "111111" when address = "0010110011101" else
            "111111" when address = "0010110011110" else
            "111111" when address = "0010110011111" else
            "111111" when address = "0010110100000" else
            "111111" when address = "0010110100001" else
            "111111" when address = "0010110100010" else
            "111111" when address = "0010110100011" else
            "111111" when address = "0010110100100" else
            "111111" when address = "0010110101000" else
            "111111" when address = "0010110101001" else
            "111111" when address = "0010110101010" else
            "111111" when address = "0010110101110" else
            "111111" when address = "0010110101111" else
            "111111" when address = "0010110110000" else
            "111111" when address = "0010110110100" else
            "111111" when address = "0010110110101" else
            "111111" when address = "0010110110110" else
            "111111" when address = "0010110111010" else
            "111111" when address = "0010110111011" else
            "111111" when address = "0010110111100" else
            "111111" when address = "0010110111101" else
            "111111" when address = "0010110111110" else
            "111111" when address = "0010110111111" else
            "111111" when address = "0010111000000" else
            "111111" when address = "0010111000001" else
            "111111" when address = "0010111000010" else
            "111111" when address = "0011000001010" else
            "111111" when address = "0011000001011" else
            "111111" when address = "0011000001100" else
            "111111" when address = "0011000010011" else
            "111111" when address = "0011000010100" else
            "111111" when address = "0011000010101" else
            "111111" when address = "0011000011001" else
            "111111" when address = "0011000011010" else
            "111111" when address = "0011000011011" else
            "111111" when address = "0011000100010" else
            "111111" when address = "0011000100011" else
            "111111" when address = "0011000100100" else
            "111111" when address = "0011000101000" else
            "111111" when address = "0011000101001" else
            "111111" when address = "0011000101010" else
            "111111" when address = "0011000110100" else
            "111111" when address = "0011000110101" else
            "111111" when address = "0011000110110" else
            "111111" when address = "0011000111010" else
            "111111" when address = "0011000111011" else
            "111111" when address = "0011000111100" else
            "111111" when address = "0011010001010" else
            "111111" when address = "0011010001011" else
            "111111" when address = "0011010001100" else
            "111111" when address = "0011010010011" else
            "111111" when address = "0011010010100" else
            "111111" when address = "0011010010101" else
            "111111" when address = "0011010011001" else
            "111111" when address = "0011010011010" else
            "111111" when address = "0011010011011" else
            "111111" when address = "0011010100010" else
            "111111" when address = "0011010100011" else
            "111111" when address = "0011010100100" else
            "111111" when address = "0011010101000" else
            "111111" when address = "0011010101001" else
            "111111" when address = "0011010101010" else
            "111111" when address = "0011010110100" else
            "111111" when address = "0011010110101" else
            "111111" when address = "0011010110110" else
            "111111" when address = "0011010111010" else
            "111111" when address = "0011010111011" else
            "111111" when address = "0011010111100" else
            "111111" when address = "0011100001010" else
            "111111" when address = "0011100001011" else
            "111111" when address = "0011100001100" else
            "111111" when address = "0011100010011" else
            "111111" when address = "0011100010100" else
            "111111" when address = "0011100010101" else
            "111111" when address = "0011100011001" else
            "111111" when address = "0011100011010" else
            "111111" when address = "0011100011011" else
            "111111" when address = "0011100100010" else
            "111111" when address = "0011100100011" else
            "111111" when address = "0011100100100" else
            "111111" when address = "0011100101000" else
            "111111" when address = "0011100101001" else
            "111111" when address = "0011100101010" else
            "111111" when address = "0011100110100" else
            "111111" when address = "0011100110101" else
            "111111" when address = "0011100110110" else
            "111111" when address = "0011100111010" else
            "111111" when address = "0011100111011" else
            "111111" when address = "0011100111100" else
            "111111" when address = "0011110001101" else
            "111111" when address = "0011110001110" else
            "111111" when address = "0011110001111" else
            "111111" when address = "0011110010000" else
            "111111" when address = "0011110010001" else
            "111111" when address = "0011110010010" else
            "111111" when address = "0011110011001" else
            "111111" when address = "0011110011010" else
            "111111" when address = "0011110011011" else
            "111111" when address = "0011110100010" else
            "111111" when address = "0011110100011" else
            "111111" when address = "0011110100100" else
            "111111" when address = "0011110101000" else
            "111111" when address = "0011110101001" else
            "111111" when address = "0011110101010" else
            "111111" when address = "0011110110100" else
            "111111" when address = "0011110110101" else
            "111111" when address = "0011110110110" else
            "111111" when address = "0011110111010" else
            "111111" when address = "0011110111011" else
            "111111" when address = "0011110111100" else
            "111111" when address = "0011110111101" else
            "111111" when address = "0011110111110" else
            "111111" when address = "0011110111111" else
            "111111" when address = "0011111000000" else
            "111111" when address = "0011111000001" else
            "111111" when address = "0011111000010" else
            "111111" when address = "0011111000011" else
            "111111" when address = "0011111000100" else
            "111111" when address = "0011111000101" else
            "111111" when address = "0100000001101" else
            "111111" when address = "0100000001110" else
            "111111" when address = "0100000001111" else
            "111111" when address = "0100000010000" else
            "111111" when address = "0100000010001" else
            "111111" when address = "0100000010010" else
            "111111" when address = "0100000011001" else
            "111111" when address = "0100000011010" else
            "111111" when address = "0100000011011" else
            "111111" when address = "0100000100010" else
            "111111" when address = "0100000100011" else
            "111111" when address = "0100000100100" else
            "111111" when address = "0100000101000" else
            "111111" when address = "0100000101001" else
            "111111" when address = "0100000101010" else
            "111111" when address = "0100000110100" else
            "111111" when address = "0100000110101" else
            "111111" when address = "0100000110110" else
            "111111" when address = "0100000111010" else
            "111111" when address = "0100000111011" else
            "111111" when address = "0100000111100" else
            "111111" when address = "0100000111101" else
            "111111" when address = "0100000111110" else
            "111111" when address = "0100000111111" else
            "111111" when address = "0100001000000" else
            "111111" when address = "0100001000001" else
            "111111" when address = "0100001000010" else
            "111111" when address = "0100001000011" else
            "111111" when address = "0100001000100" else
            "111111" when address = "0100001000101" else
            "111111" when address = "0100010001101" else
            "111111" when address = "0100010001110" else
            "111111" when address = "0100010001111" else
            "111111" when address = "0100010010000" else
            "111111" when address = "0100010010001" else
            "111111" when address = "0100010010010" else
            "111111" when address = "0100010011001" else
            "111111" when address = "0100010011010" else
            "111111" when address = "0100010011011" else
            "111111" when address = "0100010100010" else
            "111111" when address = "0100010100011" else
            "111111" when address = "0100010100100" else
            "111111" when address = "0100010101000" else
            "111111" when address = "0100010101001" else
            "111111" when address = "0100010101010" else
            "111111" when address = "0100010110100" else
            "111111" when address = "0100010110101" else
            "111111" when address = "0100010110110" else
            "111111" when address = "0100010111010" else
            "111111" when address = "0100010111011" else
            "111111" when address = "0100010111100" else
            "111111" when address = "0100010111101" else
            "111111" when address = "0100010111110" else
            "111111" when address = "0100010111111" else
            "111111" when address = "0100011000000" else
            "111111" when address = "0100011000001" else
            "111111" when address = "0100011000010" else
            "111111" when address = "0100011000011" else
            "111111" when address = "0100011000100" else
            "111111" when address = "0100011000101" else
            "111111" when address = "0101010001101" else
            "111111" when address = "0101010001110" else
            "111111" when address = "0101010001111" else
            "111111" when address = "0101010010000" else
            "111111" when address = "0101010010001" else
            "111111" when address = "0101010010010" else
            "111111" when address = "0101010011001" else
            "111111" when address = "0101010011010" else
            "111111" when address = "0101010011011" else
            "111111" when address = "0101010100101" else
            "111111" when address = "0101010100110" else
            "111111" when address = "0101010100111" else
            "111111" when address = "0101010101011" else
            "111111" when address = "0101010101100" else
            "111111" when address = "0101010101101" else
            "111111" when address = "0101010101110" else
            "111111" when address = "0101010101111" else
            "111111" when address = "0101010110000" else
            "111111" when address = "0101010110001" else
            "111111" when address = "0101010110010" else
            "111111" when address = "0101010110011" else
            "111111" when address = "0101010110100" else
            "111111" when address = "0101010110101" else
            "111111" when address = "0101010110110" else
            "111111" when address = "0101010111010" else
            "111111" when address = "0101010111011" else
            "111111" when address = "0101010111100" else
            "111111" when address = "0101010111101" else
            "111111" when address = "0101010111110" else
            "111111" when address = "0101010111111" else
            "111111" when address = "0101011000000" else
            "111111" when address = "0101011000001" else
            "111111" when address = "0101011000010" else
            "111111" when address = "0101100001101" else
            "111111" when address = "0101100001110" else
            "111111" when address = "0101100001111" else
            "111111" when address = "0101100010000" else
            "111111" when address = "0101100010001" else
            "111111" when address = "0101100010010" else
            "111111" when address = "0101100011001" else
            "111111" when address = "0101100011010" else
            "111111" when address = "0101100011011" else
            "111111" when address = "0101100100101" else
            "111111" when address = "0101100100110" else
            "111111" when address = "0101100100111" else
            "111111" when address = "0101100101011" else
            "111111" when address = "0101100101100" else
            "111111" when address = "0101100101101" else
            "111111" when address = "0101100101110" else
            "111111" when address = "0101100101111" else
            "111111" when address = "0101100110000" else
            "111111" when address = "0101100110001" else
            "111111" when address = "0101100110010" else
            "111111" when address = "0101100110011" else
            "111111" when address = "0101100110100" else
            "111111" when address = "0101100110101" else
            "111111" when address = "0101100110110" else
            "111111" when address = "0101100111010" else
            "111111" when address = "0101100111011" else
            "111111" when address = "0101100111100" else
            "111111" when address = "0101100111101" else
            "111111" when address = "0101100111110" else
            "111111" when address = "0101100111111" else
            "111111" when address = "0101101000000" else
            "111111" when address = "0101101000001" else
            "111111" when address = "0101101000010" else
            "111111" when address = "0101101000011" else
            "111111" when address = "0101110001101" else
            "111111" when address = "0101110001110" else
            "111111" when address = "0101110001111" else
            "111111" when address = "0101110010000" else
            "111111" when address = "0101110010001" else
            "111111" when address = "0101110010010" else
            "111111" when address = "0101110011001" else
            "111111" when address = "0101110011010" else
            "111111" when address = "0101110011011" else
            "111111" when address = "0101110100101" else
            "111111" when address = "0101110100110" else
            "111111" when address = "0101110100111" else
            "111111" when address = "0101110101011" else
            "111111" when address = "0101110101100" else
            "111111" when address = "0101110101101" else
            "111111" when address = "0101110101110" else
            "111111" when address = "0101110101111" else
            "111111" when address = "0101110110000" else
            "111111" when address = "0101110110001" else
            "111111" when address = "0101110110010" else
            "111111" when address = "0101110110011" else
            "111111" when address = "0101110110100" else
            "111111" when address = "0101110110101" else
            "111111" when address = "0101110110110" else
            "111111" when address = "0101110111010" else
            "111111" when address = "0101110111011" else
            "111111" when address = "0101110111100" else
            "111111" when address = "0101110111101" else
            "111111" when address = "0101110111110" else
            "111111" when address = "0101110111111" else
            "111111" when address = "0101111000000" else
            "111111" when address = "0101111000001" else
            "111111" when address = "0101111000010" else
            "111111" when address = "0101111000011" else
            "111111" when address = "0101111000100" else
            "111111" when address = "0110000001010" else
            "111111" when address = "0110000001011" else
            "111111" when address = "0110000001100" else
            "111111" when address = "0110000010011" else
            "111111" when address = "0110000010100" else
            "111111" when address = "0110000010101" else
            "111111" when address = "0110000011001" else
            "111111" when address = "0110000011010" else
            "111111" when address = "0110000011011" else
            "111111" when address = "0110000100101" else
            "111111" when address = "0110000100110" else
            "111111" when address = "0110000100111" else
            "111111" when address = "0110000101011" else
            "111111" when address = "0110000101100" else
            "111111" when address = "0110000101101" else
            "111111" when address = "0110000111010" else
            "111111" when address = "0110000111011" else
            "111111" when address = "0110000111100" else
            "111111" when address = "0110001000011" else
            "111111" when address = "0110001000100" else
            "111111" when address = "0110001000101" else
            "111111" when address = "0110010001010" else
            "111111" when address = "0110010001011" else
            "111111" when address = "0110010001100" else
            "111111" when address = "0110010010011" else
            "111111" when address = "0110010010100" else
            "111111" when address = "0110010010101" else
            "111111" when address = "0110010011001" else
            "111111" when address = "0110010011010" else
            "111111" when address = "0110010011011" else
            "111111" when address = "0110010100101" else
            "111111" when address = "0110010100110" else
            "111111" when address = "0110010100111" else
            "111111" when address = "0110010101011" else
            "111111" when address = "0110010101100" else
            "111111" when address = "0110010101101" else
            "111111" when address = "0110010111010" else
            "111111" when address = "0110010111011" else
            "111111" when address = "0110010111100" else
            "111111" when address = "0110011000011" else
            "111111" when address = "0110011000100" else
            "111111" when address = "0110011000101" else
            "111111" when address = "0110100001010" else
            "111111" when address = "0110100001011" else
            "111111" when address = "0110100001100" else
            "111111" when address = "0110100010011" else
            "111111" when address = "0110100010100" else
            "111111" when address = "0110100010101" else
            "111111" when address = "0110100011001" else
            "111111" when address = "0110100011010" else
            "111111" when address = "0110100011011" else
            "111111" when address = "0110100100101" else
            "111111" when address = "0110100100110" else
            "111111" when address = "0110100100111" else
            "111111" when address = "0110100101011" else
            "111111" when address = "0110100101100" else
            "111111" when address = "0110100101101" else
            "111111" when address = "0110100111010" else
            "111111" when address = "0110100111011" else
            "111111" when address = "0110100111100" else
            "111111" when address = "0110101000011" else
            "111111" when address = "0110101000100" else
            "111111" when address = "0110101000101" else
            "111111" when address = "0110110001010" else
            "111111" when address = "0110110001011" else
            "111111" when address = "0110110001100" else
            "111111" when address = "0110110010011" else
            "111111" when address = "0110110010100" else
            "111111" when address = "0110110010101" else
            "111111" when address = "0110110011100" else
            "111111" when address = "0110110011101" else
            "111111" when address = "0110110011110" else
            "111111" when address = "0110110100010" else
            "111111" when address = "0110110100011" else
            "111111" when address = "0110110100100" else
            "111111" when address = "0110110101011" else
            "111111" when address = "0110110101100" else
            "111111" when address = "0110110101101" else
            "111111" when address = "0110110101110" else
            "111111" when address = "0110110101111" else
            "111111" when address = "0110110110000" else
            "111111" when address = "0110110110001" else
            "111111" when address = "0110110110010" else
            "111111" when address = "0110110110011" else
            "111111" when address = "0110110111010" else
            "111111" when address = "0110110111011" else
            "111111" when address = "0110110111100" else
            "111111" when address = "0110110111101" else
            "111111" when address = "0110110111110" else
            "111111" when address = "0110110111111" else
            "111111" when address = "0110111000000" else
            "111111" when address = "0110111000001" else
            "111111" when address = "0110111000010" else
            "111111" when address = "0110111000011" else
            "111111" when address = "0110111000100" else
            "111111" when address = "0111000001010" else
            "111111" when address = "0111000001011" else
            "111111" when address = "0111000001100" else
            "111111" when address = "0111000010011" else
            "111111" when address = "0111000010100" else
            "111111" when address = "0111000010101" else
            "111111" when address = "0111000011100" else
            "111111" when address = "0111000011101" else
            "111111" when address = "0111000011110" else
            "111111" when address = "0111000100010" else
            "111111" when address = "0111000100011" else
            "111111" when address = "0111000100100" else
            "111111" when address = "0111000101011" else
            "111111" when address = "0111000101100" else
            "111111" when address = "0111000101101" else
            "111111" when address = "0111000101110" else
            "111111" when address = "0111000101111" else
            "111111" when address = "0111000110000" else
            "111111" when address = "0111000110001" else
            "111111" when address = "0111000110010" else
            "111111" when address = "0111000110011" else
            "111111" when address = "0111000111010" else
            "111111" when address = "0111000111011" else
            "111111" when address = "0111000111100" else
            "111111" when address = "0111000111101" else
            "111111" when address = "0111000111110" else
            "111111" when address = "0111000111111" else
            "111111" when address = "0111001000000" else
            "111111" when address = "0111001000001" else
            "111111" when address = "0111001000010" else
            "111111" when address = "0111001000011" else
            "111111" when address = "0111010001010" else
            "111111" when address = "0111010001011" else
            "111111" when address = "0111010001100" else
            "111111" when address = "0111010010011" else
            "111111" when address = "0111010010100" else
            "111111" when address = "0111010010101" else
            "111111" when address = "0111010011100" else
            "111111" when address = "0111010011101" else
            "111111" when address = "0111010011110" else
            "111111" when address = "0111010100010" else
            "111111" when address = "0111010100011" else
            "111111" when address = "0111010100100" else
            "111111" when address = "0111010101011" else
            "111111" when address = "0111010101100" else
            "111111" when address = "0111010101101" else
            "111111" when address = "0111010101110" else
            "111111" when address = "0111010101111" else
            "111111" when address = "0111010110000" else
            "111111" when address = "0111010110001" else
            "111111" when address = "0111010110010" else
            "111111" when address = "0111010110011" else
            "111111" when address = "0111010111010" else
            "111111" when address = "0111010111011" else
            "111111" when address = "0111010111100" else
            "111111" when address = "0111010111101" else
            "111111" when address = "0111010111110" else
            "111111" when address = "0111010111111" else
            "111111" when address = "0111011000000" else
            "111111" when address = "0111011000001" else
            "111111" when address = "0111011000010" else
            "111111" when address = "0111100001010" else
            "111111" when address = "0111100001011" else
            "111111" when address = "0111100001100" else
            "111111" when address = "0111100010011" else
            "111111" when address = "0111100010100" else
            "111111" when address = "0111100010101" else
            "111111" when address = "0111100011100" else
            "111111" when address = "0111100011101" else
            "111111" when address = "0111100011110" else
            "111111" when address = "0111100100010" else
            "111111" when address = "0111100100011" else
            "111111" when address = "0111100100100" else
            "111111" when address = "0111100101011" else
            "111111" when address = "0111100101100" else
            "111111" when address = "0111100101101" else
            "111111" when address = "0111100111010" else
            "111111" when address = "0111100111011" else
            "111111" when address = "0111100111100" else
            "111111" when address = "0111101000000" else
            "111111" when address = "0111101000001" else
            "111111" when address = "0111101000010" else
            "111111" when address = "0111110001010" else
            "111111" when address = "0111110001011" else
            "111111" when address = "0111110001100" else
            "111111" when address = "0111110010011" else
            "111111" when address = "0111110010100" else
            "111111" when address = "0111110010101" else
            "111111" when address = "0111110011100" else
            "111111" when address = "0111110011101" else
            "111111" when address = "0111110011110" else
            "111111" when address = "0111110100010" else
            "111111" when address = "0111110100011" else
            "111111" when address = "0111110100100" else
            "111111" when address = "0111110101011" else
            "111111" when address = "0111110101100" else
            "111111" when address = "0111110101101" else
            "111111" when address = "0111110111010" else
            "111111" when address = "0111110111011" else
            "111111" when address = "0111110111100" else
            "111111" when address = "0111111000001" else
            "111111" when address = "0111111000010" else
            "111111" when address = "0111111000011" else
            "111111" when address = "1000000001010" else
            "111111" when address = "1000000001011" else
            "111111" when address = "1000000001100" else
            "111111" when address = "1000000010011" else
            "111111" when address = "1000000010100" else
            "111111" when address = "1000000010101" else
            "111111" when address = "1000000011100" else
            "111111" when address = "1000000011101" else
            "111111" when address = "1000000011110" else
            "111111" when address = "1000000100010" else
            "111111" when address = "1000000100011" else
            "111111" when address = "1000000100100" else
            "111111" when address = "1000000101011" else
            "111111" when address = "1000000101100" else
            "111111" when address = "1000000101101" else
            "111111" when address = "1000000111010" else
            "111111" when address = "1000000111011" else
            "111111" when address = "1000000111100" else
            "111111" when address = "1000001000010" else
            "111111" when address = "1000001000011" else
            "111111" when address = "1000010001101" else
            "111111" when address = "1000010001110" else
            "111111" when address = "1000010001111" else
            "111111" when address = "1000010010000" else
            "111111" when address = "1000010010001" else
            "111111" when address = "1000010010010" else
            "111111" when address = "1000010011111" else
            "111111" when address = "1000010100000" else
            "111111" when address = "1000010100001" else
            "111111" when address = "1000010101011" else
            "111111" when address = "1000010101100" else
            "111111" when address = "1000010101101" else
            "111111" when address = "1000010101110" else
            "111111" when address = "1000010101111" else
            "111111" when address = "1000010110000" else
            "111111" when address = "1000010110001" else
            "111111" when address = "1000010110010" else
            "111111" when address = "1000010110011" else
            "111111" when address = "1000010110100" else
            "111111" when address = "1000010110101" else
            "111111" when address = "1000010110110" else
            "111111" when address = "1000010111010" else
            "111111" when address = "1000010111011" else
            "111111" when address = "1000010111100" else
            "111111" when address = "1000011000010" else
            "111111" when address = "1000011000011" else
            "111111" when address = "1000011000100" else
            "111111" when address = "1000011000101" else
            "111111" when address = "1000100001101" else
            "111111" when address = "1000100001110" else
            "111111" when address = "1000100001111" else
            "111111" when address = "1000100010000" else
            "111111" when address = "1000100010001" else
            "111111" when address = "1000100010010" else
            "111111" when address = "1000100011111" else
            "111111" when address = "1000100100000" else
            "111111" when address = "1000100100001" else
            "111111" when address = "1000100101011" else
            "111111" when address = "1000100101100" else
            "111111" when address = "1000100101101" else
            "111111" when address = "1000100101110" else
            "111111" when address = "1000100101111" else
            "111111" when address = "1000100110000" else
            "111111" when address = "1000100110001" else
            "111111" when address = "1000100110010" else
            "111111" when address = "1000100110011" else
            "111111" when address = "1000100110100" else
            "111111" when address = "1000100110101" else
            "111111" when address = "1000100110110" else
            "111111" when address = "1000100111010" else
            "111111" when address = "1000100111011" else
            "111111" when address = "1000100111100" else
            "111111" when address = "1000101000011" else
            "111111" when address = "1000101000100" else
            "111111" when address = "1000101000101" else
            "111111" when address = "1000110001101" else
            "111111" when address = "1000110001110" else
            "111111" when address = "1000110001111" else
            "111111" when address = "1000110010000" else
            "111111" when address = "1000110010001" else
            "111111" when address = "1000110010010" else
            "111111" when address = "1000110011111" else
            "111111" when address = "1000110100000" else
            "111111" when address = "1000110100001" else
            "111111" when address = "1000110101011" else
            "111111" when address = "1000110101100" else
            "111111" when address = "1000110101101" else
            "111111" when address = "1000110101110" else
            "111111" when address = "1000110101111" else
            "111111" when address = "1000110110000" else
            "111111" when address = "1000110110001" else
            "111111" when address = "1000110110010" else
            "111111" when address = "1000110110011" else
            "111111" when address = "1000110110100" else
            "111111" when address = "1000110110101" else
            "111111" when address = "1000110110110" else
            "111111" when address = "1000110111010" else
            "111111" when address = "1000110111011" else
            "111111" when address = "1000110111100" else
            "111111" when address = "1000111000011" else
            "111111" when address = "1000111000100" else
            "111111" when address = "1000111000101" else
            "111111" when address = "1010010010100" else
            "111111" when address = "1010010010101" else
            "111111" when address = "1010010010110" else
            "111111" when address = "1010010011001" else
            "111111" when address = "1010010011010" else
            "111111" when address = "1010010011110" else
            "111111" when address = "1010010011111" else
            "111111" when address = "1010010100010" else
            "111111" when address = "1010010100011" else
            "111111" when address = "1010010100100" else
            "111111" when address = "1010010100111" else
            "111111" when address = "1010010101000" else
            "111111" when address = "1010010101001" else
            "111111" when address = "1010010101010" else
            "111111" when address = "1010100010011" else
            "111111" when address = "1010100011000" else
            "111111" when address = "1010100011011" else
            "111111" when address = "1010100011101" else
            "111111" when address = "1010100100000" else
            "111111" when address = "1010100100010" else
            "111111" when address = "1010100100101" else
            "111111" when address = "1010100100111" else
            "111111" when address = "1010100101101" else
            "111111" when address = "1010110010100" else
            "111111" when address = "1010110010101" else
            "111111" when address = "1010110011000" else
            "111111" when address = "1010110011101" else
            "111111" when address = "1010110100000" else
            "111111" when address = "1010110100010" else
            "111111" when address = "1010110100011" else
            "111111" when address = "1010110100100" else
            "111111" when address = "1010110100111" else
            "111111" when address = "1010110101000" else
            "111111" when address = "1010110101001" else
            "111111" when address = "1011000010110" else
            "111111" when address = "1011000011000" else
            "111111" when address = "1011000011011" else
            "111111" when address = "1011000011101" else
            "111111" when address = "1011000100000" else
            "111111" when address = "1011000100010" else
            "111111" when address = "1011000100100" else
            "111111" when address = "1011000100111" else
            "111111" when address = "1011000101101" else
            "111111" when address = "1011010010011" else
            "111111" when address = "1011010010100" else
            "111111" when address = "1011010010101" else
            "111111" when address = "1011010011001" else
            "111111" when address = "1011010011010" else
            "111111" when address = "1011010011110" else
            "111111" when address = "1011010011111" else
            "111111" when address = "1011010100010" else
            "111111" when address = "1011010100101" else
            "111111" when address = "1011010100111" else
            "111111" when address = "1011010101000" else
            "111111" when address = "1011010101001" else
            "111111" when address = "1011010101010" else
                    "110000";




	end if;

	end process;
	
rgb <= rgb_signal;	
			
end;